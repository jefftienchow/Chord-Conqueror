BZh91AY&SY��4� �_�Px����������`	?x���,  ��cFR�Ih�0���=54di��@�@�S�2
�54d� F�� h*~�P F�     	4������ d��  �&L��L �0L�0�RB F�hSĘ�� 4P��	��� MD�!^����HlT	���{r�&��$6��Fi�X��׫�q?�'��=ݹKimˌR�[e����m-�Z[q�b  �B�D(UJRU(P��0��J�
Z�6�Җ��ڶ��[e��ۜu6[w	}�
��'�k�����v���Et��Z���´�1��t]\/�2�����uڌ����~M���I2���9O'E�R02壻��a�c%ƴ�Q��T�õ��ԯ��=�r'���/�ьp"�ǷHu#�&�T�-,q���7s �^մ�@&�Wva �0M��
J[�(7M��dC9\d��2$R��Y��g�<Z�N�� ���]{�@�aI$`���~��ͦ���fѥ�jH&'��Z���v%u����\o�cdi��q�HGö4@J�5����]�����wx+�y�J�O�X�ǟ�c�ȏ<�~qI�0:(	����l��nn�T�n��\���
EB��&�U�S5��qn���ɚ	�%�G�@V��:�gUu_(��Z��# �Rkk���<M�yx)�w*%u���l���qu8�*��É9~Nv���Z*��v+{�
�m�����B�H������&��.���Tt��>65���]�C���31u��Vb��d�x�i�Qz{��ݛ�9:��i)jv�7���0����>ɮ��z85ɟS�fo�;qF']&����_Z{�ӑ�S��{��aBA	+ �X-�L\NpHZf��B8�;!�3]�O#|�:qGQ���g,J	�6EmdQ��Z��Z�F]yN��p����L�غ'��X�U��T�Ӄ)�2�[�S�av�qWS1,�킝�WV,F���$D̻����P�����T�[������
FN�j���n0jZG��;�s箩2�!738��%Lhʃ�s��"���Cn��e��Q��nc�Zx��unq^�&�٭�;�M�هM�<��QE�UVH�,��o�=}�<+�U�|�»������z���"<im"E�*�ڪ^#��T��sJC,)��"B�#���r	`b���u�D0��p�P��H,�g���y�ޔ�Ĩ��\Np����f��u|�Ra�$k�	����(��ݙ�����j�}�fQ��p�i5#�qg��wG!�owޝ��q�6t�DFe�c���y����ʞ�G���a�O����*s�I<$DyF�{7�����4�:*�۝ɺM$�P��)�5���Zf�6�r;�"�9iu�h�4�v�~����(���-Q!�:�b��g��래j��S��p3��<�AJJ�$U��ۉ�<�ͼA���cE�a8NC�p��Wp02B����DDm�G@_�~�D�x�`��a�2�Ao hU�^AWaF���"��Y�q��5}Opk����$eYsH��;ޑI׹�C��cvf�a����l�F�ӆ�b�1}4��~�V��$�L�b�9d\��uﵮ��Z��[)����Q/X�������(��O����sH��׏M�����`#�o��Ptm*"#t�f��ax�)��;;�,"���D��Ru�9�Dq�3���M�-qׯ�FJ�Z���%.0����R�l��_���("ʄS�5�Q��1/Z�bDFM<�,�����KC��YRR����-r)2.�&�E���ԙ��@�[xR�1���E�s�G~��.ÁF�uV��7�U����H�
��� 