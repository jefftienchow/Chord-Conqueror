BZh91AY&SY#�/ M_�Px����߰����`
y���[>ؠ  �ރϟv��ܴH�4򞒞���bmCjPɠ�hѠJ�@$��`����L�����Q� 4dh �    JdD�e!��4�2i� @ IO(��1�l���244�##'�0�FjD��Sj �   � ���j*�D������{@�}Q�P��Ă��E��.��P�Q��������|�d�eS*�T�T�TʦU8�eʦU8�G	���J
BUl��L`���LL��*��r hDf�%B Js-J �
�
J�'Z�Y8����;b���~��*I�bIgY�h�M�5��\Ic)skM�Q��k3D���&�b�'y�a�cűQ�bl��K���6Jr'�TMaQo�Qk'eY�{#�x��-��^��RK2Ū� ��}�������7��n��I:ظ�a�I'�c�W�c�@%
ɼ9��|>�Mg����o�z1�ѱ��[wP\_/�h�h�iiZV�APe�Ye�n��n�����1��a�i��i�����4�Ba�����Ƶ�-"z���F�*UH�r��f�ZP�Br]Jv��b����1C̻<��)���%�Xy�&L���E�^�2.W#� �8��`X�X�X��L���[C|�)�����H�M�W�	�H˘ҧL��E�h�"��9�jMێj2�f��#���L��c#�x�]ݎAz8�:�%���6���H�M���8plk��!
��Z,�C/��Ƒ��&R�6�<�t�l�5�t�1b�dq��h."`�WX|��:�%�è�I9�gy�$�v~�� �z ��˕f:ãi���*��~w����y�HI&ڌ�X$�G�����9�D>�~��Awd��6�q�^�h�d�~r0nG`���h<�p���6<��_��fa�{ �M���&��[��z�M��
����7Kz��L1��Ʌw�����xv%�'P�h��I7�D4i23��N���H�F �J4UR���B6N�SЗ"H�.��VP�=(z�Wzt�c���s���t�%�;;t@��n\��'���Xw��)��BI�A�)A04�I���M�;��67���$������Y�"�Fl$f���F�̒`}"`UC�VW4�n���S4u��o���HE�2��:1P`Ĕ֤r͹#��'�}�8͕$����C<�L�	�v���vnX�q+���5g������9�*Ms5sklt!�Ul��Ck�f��(��O*��O��9��?��:lxu��t�ѻ��_-¢��ɚaOa		$&˂I��P�]ԏ+(�w��AY#Љa���\sJ�K�4������sRc;k���l�EEw�P@�*+׮��ÅR�LB�J���A͈e���D#$bDH�"q�l�K	"	"$A#1#cIAADQA@�d(D(����adX\�0�B�-(��ڨ)�3�l�Q	$ Y��s�o'C�q����]�O�<^�#��_Z�R�rc�̦��s]�3��,/��ޥi�0� .���<���^�p���K ��j�Fr���gbI$���Z�uT}�E�5��} ��p�f�����]���Y҈�|_�v�\;�Zn���.ay	rXI -G\���Jp�b9$�iA!��B%�n)k|� �ň6�s��%IRpV?vH�V$��9qX��b���N��{Aۖt"I<�<�1~��脭&�HQɘo
��Do9\3ؘ.1@���Q��8�춛ס٣�dca�n-���������H����.‘�c��ם�#8��h�������'*��{y��l�D�B�-��npOE����ѐ��,0�}1��0��S��0cc
��dC��U��ʨM�]Tڤ��,C�p�ra�&Ӣ�J�(�1��yW���N�*""�8��ojj�pQ`�jl���e�2;ނ���.�����49�7.��f]�,��q��m`dc���)���x