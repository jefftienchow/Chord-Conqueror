BZh91AY&SYD�j� G_�Px����߰����` 8 wX          `�J���� ��Ț�����I�h�i��5<@*J� 41222h!�101��&F�ISA� �     ѓ �`A��2`�$����=�=�R?T�O(4�OMji��WT'B��H��P�DP�g�y���c��
���%�E2"����^9OGA���~��>�U�Qb,��YE���(�Q�o�4,й�H�e"�,E��YE���e"�,E���,E�Y�f��hX���H3(�B�Y�b,��YE��0&	E���1Qb,��YE���e �(��YA&����YpX���f��S1Q�"�h�E����b.e�b,�� ሱQ�f��u���;�N��-�%��v����3+�,��.F$�o�Nꊩ��qF�ԡD�Ћ�ə���D�ˋ�z�S��Y(�G����f����F蝨�.D���㔊���Q�#U�*�׎�Ez��gPfg=����;��6�a�$��;�nR��w�S�N|����y�"F�AB�kU{R6.n�Vvl�1z+e� �n�Q��ܯ]�bf
��r"*�FaTZ��62��Bm�������Ff
�{�Jr�,�L���wQ���;V�Ҽ��Z�4��P�U#3*f���"QJ�e݈��16	X�Sq6L���d��gaC;���_����wRDI����G+�^ay"P�+�U �͖P@4����NM�Р(B0������kdVP/�u��6��ڶJS�'	(�:�"�jO��՜¬4��ث�a���p>"�N�t|�v����P���5�TȄj\��۴6��J��U��cF�Я�YTlM����f�L�uЄ.��$$K�����bWV(��,[��m�v#�T%�O��n�ڭ���෵��r��LQc�V���2����$�<:�� {�Dx|��Fˌ���OU9�)�BӬ���(B��m��x�����{�
{��Ǝ��CcDvA6)X��K����� q��˵�B�,IcK�`����jb2%q�0R�v1��E�P���!���k�һ����R$�C�:j��n�0���:�R�9#(:(U7R*#.!��x":�|g�@�>��J�6����1a,�I��z���|�����h�w�j��o.�Xx�����5
o~a�H(�������.���H��1N�������Ҵ6��\	�HbnVGh%��oU��<�̡J���iJ\�z��12.�ȑBT����a0��"8��y�	�;���*8bLO)�c��:ʉ,!�Xv�i��&�H'h@q�0��"8!k7�x�X��R����z笙V�Ae��v�qR.��	�S6�",V*qg$hb�]����0�\�X�GT�`��ɳ�2��V��
�"�U�oP��Ch�I�}�E��ˇS �ݘP ���sb�T#FIi��EA�F�o ���#���[��5���Q��C;th���fޜ�pCy��NN#�nԛ� r0F����r�Ŵ�7-Jb�6ౖ��ܡ�y�����0�ڬ34%H�V\�E��q�<+�����
Y�����$+�d�Vl�x�.�z}u[��$#	DFm읰)n
LC5n�UXW�#�!��5әT���dq��6!��T:硃	]�9f�n��
a��T�TXi��8_;�^2e�U1�8`A�$h�R�8^�c/5B��Ƴ�ES4)���am�<P����7�O��F�؟���8C �4X�},�aV���S��_AΥYA����ND�P/��6�I��y�4�T�Qہ�1r t���42"�ĄՌ�f!s�HU�p�
�ݸ������(sd1��;H+&�{��AV�c����c_�X�X���kH�M�5r���P����H�4a�=�f$����M`g�@���s9:bb
X�9"����q���s�Yf�mMC���l>wuJ�\R��y�T�H�C��.�)d�S��yv�K(�+B���%�LX6���д���U���9��oz���ŝ���!�,�NsCd�hT��{�5�I{7C!�)���#�Y��0cM@�������`,�����n	�@#/����G��t>�
�ЎRt�z��׈L���� 翤�B�pZ\ed��V�M���N�Kd���mR�N]�chv�DQ�j�5U+���]��ڬ��Ц���	��rPBD&�.C�qT��� ��`I�B����T���ް�Q�(�İ�c�t3��ι2w2�g����0eG�)�f>��sV�����}!�O����$L@��&1-�ṝP�g�#�	#elz�ҹ���՜J��JW�1�/(3*m�|�y�W�}|�Y�͹�;!ȯ�!hj��^����6�L���7�OD��2),l1�*a�d����!����fhߟ<��~
�z�W;3YE⋐ЁH�Sudr�J�X(��9�'�\�	
�/B�xe�ڜӻd���P�N'��DX�x2T�BP���0M����0W��8CW��I�%��F�F��u�2�Q9��	Y]�0Z$�fáb��aDn������D�#Dr�Bn�le��0�s�"���DC��2ϭE�(!��pVYQ�t��b�b��=^�a�����^�S������\���UQg�Be��\�<5a��萄���I @AB�:z�GuwqX��Am��u�������cC�ک.@%B�� ����ԑ�dX��Ҹ4Zg-����}f�zPD�G�x�k�>��r�i�WY��РZ�����$0��H���~�I��^��ϗe.�co����Ӣ��� H:������O*�w�]@P�R��uN�f��u����6s>$9��P>߻۰�.���YZ�h|&T��g�,�$;�)U\����wbШPc�e�`�!�A�P-cp�+T燨�D��5�C�c�YW�RZ��p��Y��W�#��$S��p�q�����y�w�x��q��m��ݗ`k�!�xtbX`�q r[�)�K
�	 �R�a����d��,�(TPڠ(}9�;��7���U��9Q��q^A�Ԓ� �t3 i
><�g����T�w�m�1�b�&㲙Ē$�����!�i�@P�Xwq�E}Gv}����ϋC��X�42���2;���6*D$}��'r�Ԡ(l�e����7g���ɪC4�_!dgL5�-�JLa��ʐ���t��BA[�H%Mc��9�BчFbA�]U�t����hΏ��Z��ʧ����n9:�ek2�1R�'Vk�å���[u��w$S�	Iv�