BZh91AY&SY�(Gt R߀Px������?���Pٞ�.Ŷ�n��D�&�jOS�OMM=!���F��=A��cS
L�SF���     H�"��4���Q��z�( CL�9�&& &#4���d�#�)�4F�$d� h  hh8(�$�PEĠ�����(�H:�᯼��H��Y���B����z>�|=;�l�k�M�a}��J��d��Pd��K����2a&��(xxu�.C� +��m�J�� FS@H$sf�����hա�ص�&.���2��0��K�65K.����Ԯ^Q�$P�G�ʌ�x��d��ad�1�a��*��3��H�iE�wjP���:7[cco�i�9{����-�cqBe���8R\�E�������#m1��X.��j��a���D���k�ef��0gNX<��»�Ӧ[��O3�����C�Q�F��Q�ņ�YP�tϺ�*�[?>�]o�Q�]��4�9�.���� 9�N<gn��y�G���4��~�Z<Wx���y��,c+]3�8R���`o�ȋ)][���Pau�𵑳�S�����6Ug��
��'L�yI�as|�=�>��{�2_�g�+�R��>�Z߃���	Ʊ�Z��
�PF0��<��0I�B
�ZC:ަ<���W7g܋dZ�p8v���oR�i��L�p���.CtLb�E�X"LX���'� ��a��� bQ�I��BRP�3��:�C�!�*I���b���Ne�=�W�~(t�hp��
�i��pkoL��p+��)'�N��.ae�$^�*=�̍�"��Ab��눺8(��*�<P̹�L8P�Y�|���&�����2�P=�ª�m�AK8¢dxI>�!�뇑����V�.��E�,��\��$+�C��벫��9R��E����8�a�g���]��BC<��