BZh91AY&SY��k Y_�Px����߰����`� `z��t%$��H�(�@I�tD�1$��x�L5 h   �"����IS� b�  4  hɉ�	���0 �`�0�*��� UP       �2b`b0#L1&L0D�F��h�S!�F�L��i�ӋlӀ"�� (3 �UhY��h�_��*?C�t���\H�{#P#��s���ʞD�I�%$JJH���d�Y"D��I�%$JH��)"RRD��Y,�H� i,�,�)"R@
H��)"RD��I�%%JJ��B�R$K��D��F��I R@�%0"D�Ӄ���ɮ�o?��~���\L #��x���k}�Ÿ�@j��n.N�^R%�5����JU�8Z�^$c M��26&����F`� �7#]̪�^�����X���9O2��qP�w:e=WN�"X�b�����ɍ�m�
L!����L]Л́�T��]JV*�AZ���&d���=�[RĦ��1���[��2`�eLI�hY�/t!)�fSt�t32��z؍�I�-;���@��f��j�8�.��gH���-bې��g� IP��DQL%XG?@�(ca��P@4����I�� UTQ_]�Ů��&
xqș+���LH�`CRQ�2��4��\��OdQ�搮�-��x0���88�+��B�>hM2mmN��U��d�]lk���i�[�v�4?*��K^eVbqM��2�1,�N�OT:Q�a�Vb�8���3��t4s#3n@h�
�R[b�`�n� Z8�Nz�#̳�ɽ�9+mRS
*l�GekɁ]��c��w+�a���QJn�ء��`�MX*h�TNIe�]&��3���U�s�6`L��k'��j��1�^����,sQ�=�p�j��b5s�I��5H�A3��e.X10�.�,��er�3�q�{V×s��yJ��@Kyv�j�oLt��	��F�b�8�*�{�VM���[{�huT�q��Y���4���NZ�{6m��l�Q3@;�콵A�9�1)PL�1�2
��*�.�@�[��w �A�ː*G3ػ���]}N0�]�F�
�#�L �����ֻ�9��]0�7�f���4Xr��d�.bM+���E�3v��J4�=7��D�[d�*Q��\-��3s-�q�%�Rt�A��cz�r���GOr -ۤ��a�Trp�[���R���k�b��:����ys��*H$,�v�k�o�nl�#�4L����Ծ�]��&2�� 6����b�k��J��rkq�ph���Cu8ECo2������(�6�WfT����H��̺H,�|��D4���͉3UY�lk�Tٝ�Ri;Gr�dd�l�:����DpT	ܣ�U�M	=�HdP[�Y����}J����7�D����)��9A��R�2������p�EZ�y���$�͙���^��>�51�*97���\�sz���]����0�&L&,z�3&���s�N�b��[Q�2z�l�xi ��-v�g��M9�Z�D����$޻�3��'zej�Dś�^j���gG\��\�j3�H9��;Q=ʥ�u��4F�@��C�^�Ed͝c.:T0��g�
;S�u����<[JR�PUθ�b�\d��ݫڋ��C&*�@P;`
4���0��`�]0�kr;C�ٚH�w�����vzur��rDvt�ؙHJ�e�t�{>f�E)��}W�Ɣv�0���
�쬮�R�]X���q�S�]�Cy�;����U�tQ�xOL,����(d{�#�"�td���ɖ���M�@܁w�j}���>�Ͱ�����]*9�`�b�2�y�`���$ҎQ8)�H]OO9�Qxc�B�&ƽ0U�
SU�����/U���̹�Y��ʉ-�ܛ��u��M�&�c�d�����tne���<�W�z�2��]�Q��oѹ��%GX8���d����{zz�G{Y5Χ�91��dS�]��)Y����njfj`E,��;@̎1���VV��GLo[���*�]���,��<�Fq���|�yQ2v	콫y�����8pR5|�'�V�p�nT�ί(�"�ׂ�sz�#.��7h��.�:s��e��+N���&�Gt3r:&2�����h%����4l��;\:U���|��tM�/",*F@H�u�����k��]F��9x�۹�@�g���a1���*32RTb��ܢ��z��� @�$�"�s�r�(<�b�%�*�t[Z]yik��W�٨P0�PQP- �HT��>q�nh��-���|}&[�EAD$tϕVS��^�p�1�ǣǷ���/���"����Ǿ�Dw��z����?F�����Ǐ"?��λ�۳�5�*�]Xm��޾�ǚ *ة����w�a�`�:II��9��� *���ûa�0Hn�a6��� �@�4\�޳N�D�{�2�Gf�Z�A��d/W���G�:*�T�!�Bwt��>�
���p/�+�H�ߟ�qP׉�����_{�ө� kYOIg����׸�۳R�6N�����ic��[C�~���\x�'x�'�S��]����n�J*��|�#�0xt�<����@q�B_C��i��+�p㶒�*�4B��Ƣ���E_Lj~�^N�١�!��(��v��*�pN�/xI�o �Qa���+���ߎ��.[^�&x1!a9f�!v�@R����܀�5hSCD{���v�\�/N�z�L�Ҍ��$�#t���{u����8���ǇbׅŴep���U[��D)0Q�P~aix��@�OI��$'��*B��c!Ev2vYB�|���q݂r��D̠�S?���)��_{X