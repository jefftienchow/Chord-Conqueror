BZh91AY&SY�hg #_�Px����߰����`�q�`  �)���	"L�#	45?T��M��L��h�!��)�JP ��0�M  sbh0�2d��`�i���!�i�!LP ��@�� d���&L�20�&�db``$MA2d2��i�j~� ��dhs]DI�@@ 2AS2��,��G��� �+�Ty�yA��)��b�j���᪃���$K�	���A$h!�J!C+	��)��C2�$QNݹ����͈� ����g�]{r��v�ܨUF y~�b�eFQ�x�Y�6�/ی��;���QQ8֨N2|&�U6,0����F-!�T��J�r��!wˇ��?u]�D5=Sr��r�����t��Ȣ�`簣���||omd��@�0�x5<٬��N�(�ק',�~�*+%mD�1�:b`G�b^�E�zv�=z�6Y�N�ᢀtN��*T׊�<2�{�w���z�<�&�Q��Yno��>y�<P	��9L�B�qY5e�.������\��i"�JUo��)��qW8�N��� Kɓ0��T�u�_i%��G�ɩ�\�%MWj_u.�v),;������ޚ����e�h#:��u(
N1bC5��^�����`b���@��P�$�E�ڍȡb���N)�֓pUa�YXs�;�}W���ءw��S3�]U���W �	F����y����st����nCxۚ=-�0�����E�z���}L�O�Uْ�'_e'.�;Ϯ��4�u����΋
@��E����������$jU��15�,ɶ�f����X��l���9��]�cY�Q�˨���clKN�xl]��tI��@8�{�������E���Q���fv�N᫫��"�["DL�|8��=�X�:��^�ws��8��^z~m�양���}W|��}uI�9	���g=H�Q*cFT+�7A���f[Cn��-yT/L�y���7����.��+�b�%]-D�yY'UJpR��Y\�T�� % D��7��\�ȵ�\�m�Z_"���'�Kf�%��H�AH@��dI�F�d�E��₣\�@̒f41��cy:�r�����zT�>v���ӮA��c�vw��V]����\=��*"��sh���=�wQ�g�8�PK���A��0�3���a�wo!r$�����yPIb��q啈$��J�������d�q�:UM�sF@s=�!��ZT��%�6f��#j;�鬡S|3�Ooi��� B0DdE	\��"�r�|��&��]%Cfs��A�ގ��o�c*	[J|��wS�^=�V$��0M�A}#�oĠԠn l� ���ji:�i	��'���L_w[I��T��=r����<֎ܝ'hk3ɕ�ɮ���hY���XAH!A�i@Y��YB=O��;��@b�1���3X�s� �M�q�>N�&��ʂy�n�h�M����k�qg'2+2ٰn ����̷}�p&�g2��Z#ǿz����2.�;'B��,�(r�H!�0�6����]:�֑U�WSHD(!]�$������`ãA�Įs	mLJ���0��� Wbo
��[�̵��뱙w����Y�%�`d�?���)��C8