BZh91AY&SY���- 
`_�Px����߰����`�{����:   ���'mPI"e=LLjzJcL(��z��h4b4z�*��J��&�#4�  j?T�U@   h  h �D�� 4=CF� 2  Q$��z��@   ���=S)��Q�H z@ @ ǩ@X�EYA- +mPY>;Jp�W�0L8�j�C�n�d6�d@-Sv�Ӽ��������"�A�R)����E"��R)�R�h-��)�KU�R)E�"�H�R��E"�J(UId�E"��B)��Կ���}�}E�\y�R\�0�$�Ř-2-���kGO)<�\�<4QUY�V�Q�''�Aj5M���nM֫٧�L��kLM��SQy��u;ُ��Z3SR��[�3�E��8l���e~K����q�E��Z���w��=��
T�:#���m2Rc���8��P (D��2�����YbI!0Ɇ��-���[���E���P��wt��cL�����.n�O|"&��t��|"��N�%�T�S�L���e2�	��F�XfT�]
��J�*7XB"�R���
�'�רWIJ3���q�b���2lLJVT�_c�|}�w����Xi�e
4���L5G����*�����U�q�/4a�OqD�qZ�׽ө4�2�R\D�r/.�z�f��Ϯ���:IV���39���5�^��IM�H5)��slu˅�l���1
�ⱓ;��&qt�9�D>�~�Qݗu�XN��^�Q̱ABm��(!��[���W��\,�}^5a<Hu�jz�`沺E�ɗ�++0�"d��Fۤ(�{âSsI@��Q$޳i�$��I�;P�ɧm�[*(vI�4Uiz�j�ћȘO�Cж^��Bg��kwvc��y�k��q��CJ��ۢ��u�8h�aCߝ�R)u
�a��	�M)!�6�����-��9��Q$TX)�rDQ�,$J�ߋ4�2I�􉁪��l�4�]��T�s��D=Ty�v�S�%%+i��H�q&{���`���G�p���O"&�N	�v���z$���*��ى��>Yl�ql�<�!��.0CJ�ϯ���d�P�'�>�+�H���8�*��ey�n����*!�k�4'(��r���.���Ӯ���A�#�ġRO�er�F�ҫ�y�� Z$ݦ�PR6ߠ����B{m� �4ܻ���T���,�eҤ���/�� �a���h�#$�UJBR��A!>`$���shj�yy���Ā2g�#[����(�	d����SЗ]��	p��P%J��6%4]�kÆ=Һы??� ��9�0 �W�>ն��ߎ��d*�FVCa��0F�Ɓ��IOR��xƄ/2I!է�fP��
�v8؂(vm��^��0H)Ju��ѯ�]�����B@- #&�Bk\U��e�G۪bP���LM$��a�%��^�p<�ƃ��Fr�����#�Vޘ$����z���b·��`���m�	'��A�3��D0�M$��s0ܫ��!��a�2`��BTI$.��N�ǲ�)�-2�
�趪��.	J��dH�$�@S���%w`������@1X)�:�5Ih!�
��P"�.�E���Q�(7�v�?���C���F�q�Y���m�� c��Y��J�&����r��$����/R���z+�*٩a�(g&)6��
{�Rxf��7G6A�
��eI$�[�DDbrdd�P�n���r�eJ!���,���;��{��b3YK܋)���ٗyE�;k5�\�������"�(H{a�