BZh91AY&SY���? 		߀Px����������`	_;�   0bH$�D� "�����Q��h !�M�MF��� h4   �&L��L �0L�0�S�R�OS  �      8ɓ&# &L �# C �!���l�OI螣  OH���z(4 �a@��	�~'�c��bH��Qy��+���������D��D�ݲto���{�*�W �@P&� $�� ƢQF��n(�r���H�(� �`  �7�i�r;�=��T����ݏ�V�nӶ�&���gݑ�&�횩U7�T��W�j�`Mۋ��[^]�HSf6��i��jX��b�-vieM޵h�T��l��[�7l?��=�����=��eA���	o*�$��O�kFx�gj��Aj��j%$Z4MWD�Ü�I%UD�h�I�%e���/y-r�TH"���5c���_^fOZ���	6��?O`hȨ��+�/�_L#�����fѩ��5D��=�!���!l�v3��q��T��c�MJ����sO�*+f�vnn0m��]�Q�N칀�D�3��<�"8y�W�K\��$z��&4L )X�F}K׻�=`�U6X370.�o�xTM�{�z��K�������.߇�z�Ft�M����J��<��(���*��]yxe�[�����n�EC����@�T���= �"�,�v���:fnk��ka2a�uT�'�nD�2�"��)��;n��B�'t�5��giO_o�3�*�$;�\�0��B�x��j�qz����(`חB��-��j�����\TU���^�=ƖzXv����kn%@��.��Gl��Q]n�Z�������΋..m�(#j��p��a[6�ZX��++A�@O`�̀'V�gZ�[7>��x�%��3��+79�_vS�z�F\�5�i���M���K���X�U|�gC�`�do95L����#1CT��rw @��N�)��\����2� |jjD��,���*�{�?���� ����U��a^���Gޫ瓘|��!F� z��b4��ՕRZ-�Wve&v�.�[�z�W���eVN�N�T�w�F�;V�L���hW����� @� @$�H�ID9������xN�L�`���Z-l�Z�|����'�+<��3�[:��&/V`�r�������I�����$�R@�4@<aip�!jV��ADG�u�T$f�=�h�����?!L�KvG(@����wz���P�a�$k�	��x���dC�Ө��m`Ŭ��~��gs,j���HGP_>[V�fo���s���x9Ȣ&AHPw�a�<�.�Q��!a(c�k���
�(��M����[i�49����~�ȃ�L���{L�7��ch� ��C�'��*�&�#���1 @:A�B�:D����*m7F�I]$=�f�'LO��a2d��z�2D�1������1�Ĥ�\h2-��?}����%E=��&utQ�f@ߌ�KO,\~<s&V�-��v٘K�Q��/��!�L��pp~`�삱��<�Co@D�;"���ڢ'���O ��gl�&A���f{�ȡ6$Kܽ�N ��Kp�C����q
<m	`��ki�K�QQ>Ұ�H[eG1���2�D�<�D�������ܛTB8�#s��h��B0�o��A��H�8���j	��m���Lvl6�$����;z��=>m�"q��,����$��p�I�@�V$,B5)(�]S��!�e���S[!V�(�A���s$!)�:w2,+
�AaҜ�TTUT09\�Rd_�M�d��U�2;[���]�T�2��G��8l�n��������3��k��"��+J��H�
���