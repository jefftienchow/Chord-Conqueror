BZh91AY&SY� h߀Px����߰����`<8l�  ]q��&�K�E h!�S�z�Q�4��i������i���E?@�P�0�h a@ �0`��`ѐ��&��SjH�H����   h s F	�0M`�L"���ML�OԘ�M2  �M�UDH�PP T̪$�>��C� Y
�*	��~+�K�S8W���sn�{��8��TV��*+J��(����Ң�XYrY���%�����h�����(�����Ң��b���sr�9g�������j}���H�n�Q��T����@�X�+̅�n0&���x-�.�$)�EX4�D�,S[�J�4��
���Z�^�sE�e�Sv��s�}8Wݏ�}��Vs�&r7$�F%L,��`�E"�M+r���6�*+(��Z$��9��`%TbK��D� ��R$��߾[('5��i�G�Z��I��4���{w-��i��^W��7��u��Mf�X�v�=ztS�Q�Y5)m�0[�2J��A��ٻ�uR�pϯ"'v\�\�A��W��yyn�����D����
�T#=/�͞�w��,��]7Ł<*&�=սPE`��on<�<����޼�i�+�ґzy�(���*��\�U�o��)>�[��6��9�RZ��Ȋ����"0�3�f滰ќF�0s&���;1�l�;|�#8J���T'8�NN,��땝�={���p�D�"�'�r�T��A<a�՚���o7EJ1�з4��cl���xS����U{+��������:/�[q*>�t+������ݥ6Ǐͽ����ݤ��EU7F�gͺ�'&Lr��T�'p��i�RqWxws9�p����J��{Wݔ��ї15�i���M��].;)c]U���t;�F�}T�O��R35Kmw'r
@m���͕ˌ
1*.� ����6;v'&��,���]�[����^z�6�
�6���?R��M�]"�"�P�@��F��Z�VUIw*�n��)3�qw���7�5y��FUd���UOTw�F�;V�L���hW���G� Ԓ@�QB&����C��r%�pv'�w1�HDie�!��sX"�D���I%�� j� bU"�~%]C*t����k��D$��,g����Þ3��і�K���Jy9:���1��^H<<Yuܻ�c�+2Aj��K4-�Y��b�!�܍(N��%YY���l�S^��r�))�k�� �B�I?����'C0b�rc�h'D-�m�5��1*���^}C�t��^|�%������,TFd�a�l�c(.Ο����4	�)����CN�X�yf��*�ZS�j{+�K
�N�^2�5g�en�ۧL"�Au8����Hm$4���q5�T\�S#c�r��2�s�b�ƘV`�	7��wA���N<�a�ky�13d����kZ������k�Q /�Bν�@��G(Bh�;�9��^T��]��VR�9j��#o���H�ג���n.��z$���GS(�<J�th���g���ǁ��"E��k$;;�*	���aU*5FU"f����pLt���S35��X�@��3�v73Y���R��UA,�"fg^� ��SA`o��p[��6HO��^�u�9B���Sܩ3��瞶�q������\L
�G!w$S�	��