BZh91AY&SY�� 		_�Px����������`	?��n   nN!Q"��S ��jO�O�A�6�њF�hdzjO��*Q@��@� �  �&L��L �0L�0�M(������   �� 8ɓ&# &L �# C �!54Q�6�z��C�� 4 �h� RqE�(�E)Bi�X���� ��D�G�x^IC��T�Et�y��i"�A�v�w�c��6ص�m�����m-��Kh֖�a/	0I��� ��1110�)$�D���1.)m)im-�m-��[Km��O@uvmö_�*�7���[�w.�٧K�K� e��A�8��v�5h�J��0
�����[V�n�^ׂ���B@қ1��Pu�M�KPr�5��k�K(��n��E�4^�[�7l?��=�6������eA��*d��r��(�-#y{E�J�j7�
�Z�NBH�������pI%UD�h�E�(7O�2�g+���AD�Q��#���Ý��3~Bb�����5dXV�˱�E��\e��w'Zr��i��G�ݢ�`|�t������o�GA�95�R����sO�*+f�vnn0m��]�Q�N칀�D�3��<�8By�y�~��� �I#�zȘ�0��b��z�sg���a���M�`O
���uoTE`]O7�G�AN���>gL��M=����Ϛ��aN�b��sҦ���2�-��R}r�{���nhr [*KBډ��e�3��/e�3s]�h�#[�9�˪��8vcr$ِv�Gm��N۪����ŝ1��n�Y�Sב�f'�H.s9�aS����՚��wy�.P��.���[`�eUYs"ł��K�=ƖzXv���kn%@��.�����Q]n�Z�������΋..m�(#j��p���ٷB�ɓ���=	���8��jyl��ws9�p����D���}�O1�]s�����6��].;)c]U���t;�FF�ÓT�O��Q#1CT��rw @��N�)��\����2� |jjXiݖ9�=0���>߿}e���f�U^��U��a^�M�;<��W�&Ǟ�B�"�P�@��HՎ잫���oj��)3�qvrߍ����t#*�t�w*��c�j4�ڵ:g��KB��_} "��U�h����:����u���ܝղ���W�h��L0��R(f-�H��]�Lʼ(q-	�,P�FD0ȪXk@�3 �`b���uТg���$0�`����I��S�W��Wӫ3� z� �ٗW���H��[���nd�i����̶x���*U9�VFe����¬��a�w���4o@�o!�:�>�iv���(1�xZ�W�cv���!�E�wr����1C��}�'WB�2|(��˭�AXƛ4�:����*�&�C���1
TD�@;��R�9	A��)���v�r!������Jb�>���cǬ��O-c"f*"p��W!~�� `d�!�G\�+���⯴1ЁוI�6�HY8�<�"�P]dA�x[�S�W�0��!����pp}����`��]X-݁�bc�DO����=�'l��u����z�y\ȌH�1N��+R�*A�(,r�hK�=�[]�,U�V�j�Q� 6��ކL�d=QD����{��ξJ"{����Ľ\#4�w�t��;x$#�Nm
u�na��L}x�K�BdA!C�[�yw�(��0Gq��h���5�� MV��X�jRQ5vΎ��!ß���O�5�[���l��n먉�gYE5Fe���0:I�Х����%ܒL�;H�"��m�&G�v8�0���%35��Atj����e�:����9�����T���.�p� #-&